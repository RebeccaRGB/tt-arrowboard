/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_rebeccargb_arrow_board (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  reg [1:0] phase;
  wire [3:0] pattern = ui_in[3:0];
  wire flashing = ui_in[4];
  wire sequential = ui_in[5];
  wire lt = ui_in[6];
  wire bi = 1'b1;
  wire al = ui_in[7];
  wire [15:0] lamps;

  arrow_board ab(
    .phase(phase),
    .pattern(pattern),
    .flashing(flashing),
    .sequential(sequential),
    .lt(lt), .bi(bi), .al(al),
    .lamps(lamps)
  );

  always @(posedge clk) begin
    if (~rst_n) begin
      phase <= 0;
    end else begin
      phase <= phase + 1;
    end
  end

  // All output pins must be assigned. If not used, assign to 0.
  assign uo_out  = lamps[7:0];
  assign uio_out = lamps[15:8];
  assign uio_oe  = 8'hFF;

  // List all unused inputs to prevent warnings
  wire _unused = &{ena, uio_in, 1'b0};

endmodule
